
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CODEVHDL IS PORT(

	CLK: IN STD_LOGIC;
	
	OUTW : OUT STD_LOGIC
);	
END CODEVHDL;

ARCHITECTURE Behavioral OF CODEVHDL IS --1MHZ
	
	CONSTANT MARKSEC : STD_LOGIC_VECTOR(7 DOWNTO 0) :=X"A0"; --160 DC CYCLES
	SIGNAL COUNTSEC : STD_LOGIC_VECTOR(7 DOWNTO 0) :=X"00";
	
	CONSTANT MARKDC : STD_LOGIC_VECTOR(15 DOWNTO 0) := X"186A";		--6250
	SIGNAL COUNTER_ONE : STD_LOGIC_VECTOR(15 DOWNTO 0) := X"0000";
	SIGNAL COUNTSDC : STD_LOGIC_VECTOR(1 DOWNTO 0):="00";
		
	SIGNAL CLKDC : STD_LOGIC := '1';
	
	SIGNAL TMP : STD_LOGIC := '1';
	
	SIGNAL COUNT15 : STD_LOGIC_VECTOR(7 DOWNTO 0) := X"00";
	CONSTANT MARK15 : STD_LOGIC_VECTOR(7 DOWNTO 0) := X"3B"; --59
	
	SIGNAL FLAG :STD_LOGIC := '1';					
	
BEGIN 
	PERIOD_DIVISOR: PROCESS(CLK) BEGIN   
		 		 
		IF(CLK'EVENT AND CLK = '1') THEN		
			
			COUNTER_ONE <= COUNTER_ONE + 1;
			
			IF(COUNTER_ONE >= MARKDC) THEN
				COUNTER_ONE <= X"0000";
				CLKDC <= NOT(CLKDC);
			END IF; 
														
		END IF;				
		
	END PROCESS;
			
	DC_DIVISOR : PROCESS(CLKDC, CLK) BEGIN
		
		IF CLKDC'EVENT THEN
			IF FLAG = '1' THEN
				CASE COUNTSDC IS		
					WHEN  "00"  =>
						TMP <= '1';
					WHEN OTHERS => 
						TMP <= '0';
					END CASE;		
					
					COUNTSDC <= COUNTSDC + 1;	
					COUNT15 <= COUNT15 + 1; 
			ELSE
				TMP <= '0';						
			END IF;		

			IF COUNT15 >= MARK15 THEN
				COUNT15 <= X"00";
				COUNTSDC <= "00";		
				FLAG <= '0';
			END IF;		
					
			IF FLAG = '0' THEN
				IF(COUNTSEC = MARKSEC) THEN
					COUNTSEC <= X"00";
					FLAG <= '1';
				END IF;
				
				COUNTSEC <= COUNTSEC + 1;				
			END IF;
		 
		END IF;
																
	END PROCESS;
				
	OUTW <= TMP WHEN TMP = '1' ELSE '0';
	
END Behavioral;

